module top_module( input in, output out );
	assign out = ~in;
    // Alternative implementation
    // assign out = !in;
endmodule